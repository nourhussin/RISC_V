module cache_control(
    input wire hit, read_ready, finished_wirting,

    output wire fill, WE, RE
);

endmodule